library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package aesTest_GRBC_s18 is
  type test is record
    key      : std_logic_vector(0 to 127);
    plain    : std_logic_vector(0 to 127);
    expected : std_logic_vector(0 to 127);
  end record test;
  type testArray is array (natural range <>) of test;
  constant tests : testarray := (
    (X"000102030405060708090A0B0C0D0E0F", X"00112233445566778899AABBCCDDEEFF", X"95AF724BFB5FC72DB14642D6257ED706"),
    (X"00000000000000000000000000000000", X"F34481EC3CC627BACD5DC3FB08F273E6", X"557203D61C387E397BCD59DBFF226FD5"),
    (X"00000000000000000000000000000000", X"9798C4640BAD75C7C3227DB910174E72", X"328999B41E5FA58FDFBF8A85CA65438A"),
    (X"00000000000000000000000000000000", X"96AB5C2FF612D9DFAAE8C31F30C42168", X"B2D32D02D67BDF6F400DA6B8E0406E19"),
    (X"00000000000000000000000000000000", X"6A118A874519E64E9963798A503F1D35", X"A2AACCD6A095EC7D20565F35325FB455"),
    (X"00000000000000000000000000000000", X"CB9FCEEC81286CA3E989BD979B0CB284", X"D86C3092973B0E8542F744416B807031"),
    (X"00000000000000000000000000000000", X"B26AEB1874E47CA8358FF22378F09144", X"2016DAC838B6D84540E8D9C104659602"),
    (X"00000000000000000000000000000000", X"58C8E00B2631686D54EAB84B91F0ACA1", X"B77CE81A266B87E7617811F4CA379D9F"),
    (X"10A58869D74BE5A374CF867CFB473859", X"00000000000000000000000000000000", X"1FA5CCFE183114CB51DC2E13665BD1CC"),
    (X"CAEA65CDBB75E9169ECD22EBE6E54675", X"00000000000000000000000000000000", X"2F8BCB0CE8BEEE5C7090FF5C49678F3C"),
    (X"A2E2FA9BAF7D20822CA9F0542F764A41", X"00000000000000000000000000000000", X"BAA2D3ABD7FFDFF752B48469994BBA3A"),
    (X"B6364AC4E1DE1E285EAF144A2415F7A0", X"00000000000000000000000000000000", X"5980ED8407C70C2822D94F88915C66A4"),
    (X"64CF9C7ABC50B888AF65F49D521944B2", X"00000000000000000000000000000000", X"9ACE3A3B76907027D5D0A2CAE28B5D9C"),
    (X"47D6742EEFCC0465DC96355E851B64D9", X"00000000000000000000000000000000", X"26666663C85AD8818F43EAFE637BE861"),
    (X"3EB39790678C56BEE34BBCDECCF6CDB5", X"00000000000000000000000000000000", X"FEFF92721BE44CAF8ABC923957BD3EEF"),
    (X"64110A924F0743D500CCADAE72C13427", X"00000000000000000000000000000000", X"897DC40FF06599DC8D7D9E1004D3DE70"),
    (X"18D8126516F8A12AB1A36D9F04D68E51", X"00000000000000000000000000000000", X"5E02EC09B54847493DDECEECD2CA31D2"),
    (X"F530357968578480B398A3C251CD1093", X"00000000000000000000000000000000", X"91FBFDC0FE65AC03E07F58A57DF8AA36"),
    (X"DA84367F325D42D601B4326964802E8E", X"00000000000000000000000000000000", X"77894C6368F3ACB58B7A5FBD6C3B0CFF"),
    (X"E37B1C6AA2846F6FDB413F238B089F23", X"00000000000000000000000000000000", X"433587618979A70D61EDB4ECE5768A02"),
    (X"6C002B682483E0CABCC731C253BE5674", X"00000000000000000000000000000000", X"0E4B89ABB93DD4684EFDEC340B254E21"),
    (X"143AE8ED6555ABA96110AB58893A8AE1", X"00000000000000000000000000000000", X"79C9BC8A62843199B59AB37E7B45361A"),
    (X"B69418A85332240DC82492353956AE0C", X"00000000000000000000000000000000", X"A9713742CC55365D7DBC030779065B38"),
    (X"71B5C08A1993E1362E4D0CE9B22B78D5", X"00000000000000000000000000000000", X"C21BE1D7A488CDEAD578D84345E764D1"),
    (X"E234CDCA2606B81F29408D5F6DA21206", X"00000000000000000000000000000000", X"C86FB9FA415F626972A14CFB2A4585B1"),
    (X"13237C49074A3DA078DC1D828BB78C6F", X"00000000000000000000000000000000", X"6EBF91C1E9DA543C38F0FBD72C0BAF2C"),
    (X"3071A2A48FE6CBD04F1A129098E308F8", X"00000000000000000000000000000000", X"2B3D6A73EE6C5E2D0FB4256DB6466B6B"),
    (X"90F42EC0F68385F2FFC5DFC03A654DCE", X"00000000000000000000000000000000", X"A2DFB4B858317172B1BAA107E9B240FC"),
    (X"FEBD9A24D8B65C1C787D50A4ED3619A9", X"00000000000000000000000000000000", X"8ED156B7B9811C03B1F2492DF75BD0D0"),
    (X"00000000000000000000000000000000", X"80000000000000000000000000000000", X"18F7465093225FEB828EDEFB35C70476"),
    (X"00000000000000000000000000000000", X"C0000000000000000000000000000000", X"97563758F0CE1A744DEAEFD4351EE309"),
    (X"00000000000000000000000000000000", X"E0000000000000000000000000000000", X"20C1157697E2988EDF423751C4138BC6"),
    (X"00000000000000000000000000000000", X"F0000000000000000000000000000000", X"60874D87628389B11F5340E5F27F9F4E"),
    (X"00000000000000000000000000000000", X"F8000000000000000000000000000000", X"3F7DB90B330805D66CBE20B314771574"),
    (X"00000000000000000000000000000000", X"FC000000000000000000000000000000", X"D5CBCB441A1A77C619BF35CFE6D445D6"),
    (X"00000000000000000000000000000000", X"FE000000000000000000000000000000", X"B3691A927ED04386F82D25E2FE4E425A"),
    (X"00000000000000000000000000000000", X"FF000000000000000000000000000000", X"A66B8DF57B3C92F62968A042E36A654C"),
    (X"00000000000000000000000000000000", X"FF800000000000000000000000000000", X"25437C09A9521C0629DE8BCBC2A5AF84"),
    (X"00000000000000000000000000000000", X"FFC00000000000000000000000000000", X"1FEB9CF0F3380BF28BFDFF47451A816A"),
    (X"00000000000000000000000000000000", X"FFE00000000000000000000000000000", X"39AE71936D405DF6F59459B833564132"),
    (X"00000000000000000000000000000000", X"FFF00000000000000000000000000000", X"F8AC07E7A94EE036E44DB46F624AB151"),
    (X"00000000000000000000000000000000", X"FFF80000000000000000000000000000", X"A1B582F4E9628D2AC746DB18B7EA63B7"),
    (X"00000000000000000000000000000000", X"FFFC0000000000000000000000000000", X"2EC13DDF1ADFCD423482324A589E6224"),
    (X"00000000000000000000000000000000", X"FFFE0000000000000000000000000000", X"BE0D8CC0952C5DEC181C62F4ED54D0FD"),
    (X"00000000000000000000000000000000", X"FFFF0000000000000000000000000000", X"E34BEA8D2209AA3F6DF6E1F580297278"),
    (X"00000000000000000000000000000000", X"FFFF8000000000000000000000000000", X"0A99B5F7914DF52B38F42D98D5EC9F43"),
    (X"00000000000000000000000000000000", X"FFFFC000000000000000000000000000", X"383F0AC802C10BD83AB22593E716A1DB"),
    (X"00000000000000000000000000000000", X"FFFFE000000000000000000000000000", X"6F4A82723774A1387C77BCD8028ABFE7"),
    (X"00000000000000000000000000000000", X"FFFFF000000000000000000000000000", X"5528CA887EEB6FEADA66483467EC8391"),
    (X"00000000000000000000000000000000", X"FFFFF800000000000000000000000000", X"363B69C0661A72AC870C3559DAFF1FFD"),
    (X"00000000000000000000000000000000", X"FFFFFC00000000000000000000000000", X"A1C7944CF5D9B8B85B11E243F713904D"),
    (X"00000000000000000000000000000000", X"FFFFFE00000000000000000000000000", X"CE8FB438E42F6895A5C571258B98CC69"),
    (X"00000000000000000000000000000000", X"FFFFFF00000000000000000000000000", X"D3963D44141621380F5CDD9AAC76D4C2"),
    (X"00000000000000000000000000000000", X"FFFFFF80000000000000000000000000", X"AC1286270E0EEC9CE6D1582CEC06DC1A"),
    (X"00000000000000000000000000000000", X"FFFFFFC0000000000000000000000000", X"98076C36C149C4E06C5C226AE9755957"),
    (X"00000000000000000000000000000000", X"FFFFFFE0000000000000000000000000", X"98A8BCE1E9D100763AF3D80F2BFB520A"),
    (X"00000000000000000000000000000000", X"FFFFFFF0000000000000000000000000", X"38ACAA194641F2618FE1D62D89E62644"),
    (X"00000000000000000000000000000000", X"FFFFFFF8000000000000000000000000", X"2ED25D17AAF6F5A408AF02D8CE4A2E8F"),
    (X"00000000000000000000000000000000", X"FFFFFFFC000000000000000000000000", X"4525768D358997CF8A156F474B9F7EAA"),
    (X"00000000000000000000000000000000", X"FFFFFFFE000000000000000000000000", X"226CA220D7DE685A4588C3EB17BAC7C3"),
    (X"00000000000000000000000000000000", X"FFFFFFFF000000000000000000000000", X"DACA8E5BCEE499D908AE1F351508C4AA"),
    (X"00000000000000000000000000000000", X"FFFFFFFF800000000000000000000000", X"0072728C5BCE97BFCD84FACBDE5A1FFB"),
    (X"00000000000000000000000000000000", X"FFFFFFFFC00000000000000000000000", X"FCEB97BDFD8E71A01ECA3037C4AA4F8C"),
    (X"00000000000000000000000000000000", X"FFFFFFFFE00000000000000000000000", X"0346F6DEA24517C4C41D2028EEB5E8B9"),
    (X"00000000000000000000000000000000", X"FFFFFFFFF00000000000000000000000", X"5F1C6CE61C337B9C07221723EAD58009"),
    (X"00000000000000000000000000000000", X"FFFFFFFFF80000000000000000000000", X"AB3D937D58A6BA0D4773E46FEB9B15AF"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFC0000000000000000000000", X"5E0E35705791D4B2D4D06A11C83530D2"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFE0000000000000000000000", X"7AC8C4822351F1EB836E828554BC56F6"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFF0000000000000000000000", X"7FCF6CE4DAD494A6A2CE0D010BCF60B1"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFF8000000000000000000000", X"956A7A40FBBD30FD3CD8F5CA1D5C4C3E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFC000000000000000000000", X"1756FA3FAB849A69F8F145321C29E2C1"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFE000000000000000000000", X"BE67D64978E065A3F13B90C29C5C0AC7"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFF000000000000000000000", X"3FA08780ED7595E20EDFE438F303E24D"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFF800000000000000000000", X"3AF99CF50F70CF0CCF61E9D2D9D04DFD"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFC00000000000000000000", X"187E62B290CAEF719E2B99BB7BF5611F"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFE00000000000000000000", X"C1DB643CF38A128B7607A40646DE9440"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFF00000000000000000000", X"01BC354824A82BF0F58CDA81335B7185"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFF80000000000000000000", X"E0EB0F7CDDA52A2F62C633AF6054167E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFC0000000000000000000", X"F7238C0B2800DD68A41A31689FE50CFE"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFE0000000000000000000", X"7269C46ABED9D556B49ACCF9A92F7F50"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFF0000000000000000000", X"BA78AF77FADAA079D2A1494B96CF8DF8"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFF8000000000000000000", X"FBABCBE5BA492380122A8D3BE0C4069B"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFC000000000000000000", X"1368A3F6F9209517AE1AFE789D8F54B4"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFE000000000000000000", X"5246800249EC47E3218464FF3C4EB173"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFF000000000000000000", X"29C9C32A9E4F5DA9D6B1A9B1EB289D0B"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFF800000000000000000", X"9DD53AABE9B73A011062000BC1485C3D"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFC00000000000000000", X"80AEA8D20B9B88A25913EA1E3836804F"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFE00000000000000000", X"B9945612FA34275B182D31959DBA1992"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFF00000000000000000", X"79CB5B280FDFC99E498D7A485A83C9E5"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFF80000000000000000", X"ABFBDD9B491006E2A30C5FC336E2595B"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFC0000000000000000", X"3BABB3F159788FFF16E688132CBAACC7"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFE0000000000000000", X"820B6DBBF82F09A908F1537A2B559BBE"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFF0000000000000000", X"87610FC7A5DA98E8C3234411BD1D1D73"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFF8000000000000000", X"EB85595021D1D34C75EE287765E24A3C"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFC000000000000000", X"1C72B351837934965A0077EA82E7D4BD"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFE000000000000000", X"AA023984366C2FBF3632CA3EFA62F283"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFF000000000000000", X"5D2D57E1432B5EFD42B8A1C3364936A4"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFF800000000000000", X"F783D74F6E0B9BE1D5B68463BAF02580"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFC00000000000000", X"A530859A17B6832664DE4B5E34C14D54"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFE00000000000000", X"33E48D3590456392A00D46937AD72AA1"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFF00000000000000", X"1025B7777384A473E8761DF86B1E49B7"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFF80000000000000", X"7BD9B511D645BB07EA15F1A7A69712FE"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFC0000000000000", X"9EF7614BF20EE561F359DD8BED0B39D4"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFE0000000000000", X"BAECC17D5E85176810274654CE755BDA"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFF0000000000000", X"C6BA914199E5FE5C48587B88A7D22AD7"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFF8000000000000", X"3D049751A531F30A1E44A2ABDEA91B8E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFC000000000000", X"91AE0B55CCBC49784B2A2D9F5AAC88D5"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFE000000000000", X"DC594D9DB182EF6C6D541DC07828660E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFF000000000000", X"1BE9B7258E96E4FF6F0313237A38CF42"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFF800000000000", X"DEE73B1D39622E1248EC008079726B2C"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFC00000000000", X"8AB6A7DC6BD822BE1EC1973FBBC4C038"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFE00000000000", X"4D2766816B63D93DAC417CA65748FA11"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFF00000000000", X"132A6CF85DC85809A327E037289D1046"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFF80000000000", X"79B641245EEA656B727A8954A5564092"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFC0000000000", X"B982EBBF05FF796F5A013D5CD1FB5B70"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFE0000000000", X"C9E8C4332486AE269A190290B9ABC7AF"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFF0000000000", X"446A83ED4498582D09F1BEACE53D80CC"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFF8000000000", X"BA559B7D6F0996CA657203D3903CA637"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFC000000000", X"5987DAC0E566931A5B15C6B38C7B7695"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFE000000000", X"E5E68638BE21AD13DCDCB5BCBE99006B"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFF000000000", X"B25228E0037E4AA038688954ADBE8F65"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFF800000000", X"09F1A071F1E0E8F42C93A544C7DE739F"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFC00000000", X"9A26EA7C04170ABA4ECA9880BD90F002"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFE00000000", X"7EECA3509D402F6EAC6F14DE5A1AFF6F"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFF00000000", X"5205D94B31595854D6F24B7C11B48972"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFF80000000", X"08F04198867D95335798200168AA4AF1"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000", X"E514797BC20C5086331619A3D234BE93"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000", X"7DD5786CCF8BAFEFDC9B0A9DCC9F5047"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000", X"554DD3C1868011A359E21826890E807E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000", X"3AE06FE0CB2AB853E46AD08D9C872F78"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000", X"3656C256AA9AD8DAA224F80C912A8EC5"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000", X"BF355B267B044E3CC1D875CBC6218B0E"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000", X"66E73FB60BAEED018836AB5075FF864D"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000", X"5C5784A402D77C64698EE763A8014CF2"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000", X"7BE0F0FAC198201DEB86EB8756711090"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000", X"68E16F38DD8457B659DA239AF6F12E98"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000", X"11914C5715CF6D712B56B6CC8D9058A2"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000", X"6EF7A8962B36FD4EB6205933D8665DD3"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000", X"169CA7BF7B26AB1DFF1EFC779D0F8E27"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000", X"E70923CD743ACC883058FCF54E1D646A"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000", X"21C1CCD53A587E63DAB827D0E3BD20FF"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000", X"160ED40CCFF6D3FDC02D43FADF8387D0"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000", X"268B1F2532359C026C76E7C2F91D6871"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000", X"BB26569C4357C0A105241904C8378234"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000", X"8687945ED13D5DD6D858B7C6E26322BC"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800", X"66E9928A7D7ECA981B56D054EE566D9D"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00", X"9B5CAB8EA32709623D5297243C2A5344"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00", X"9EFBD8C3A62FD8F5A51E32E43DD4A8BE"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00", X"B1B120F3BA8BB75C241873AC54C9DAF2"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80", X"5A2F9EDA9DDFC1274EABADF0BF9A92DC"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0", X"5F5AC67F3E9A71918045AF237CF13993"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0", X"8ED195731E1C52684559F4D6A47C7B24"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0", X"61335DCD383B0094B2C4210CB2666CB9"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8", X"FDD752AF69FAD86676E5D5F1FEA29B73"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC", X"B1DB86B4179474CDFCC4900CF6592659"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE", X"877A5A8E4EE84F903AC3A8CD170555B1"),
    (X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF", X"484898A4B2B00969672968F9E1C2BC95"),
    (X"80000000000000000000000000000000", X"00000000000000000000000000000000", X"424F23300C1C68ECFD5EC70F2ABB0B93"),
    (X"C0000000000000000000000000000000", X"00000000000000000000000000000000", X"C1FF68EA3AD9AC79268268CA2F3321A3"),
    (X"E0000000000000000000000000000000", X"00000000000000000000000000000000", X"AB63AC40C4C435BF85EE75E06B8586F9"),
    (X"F0000000000000000000000000000000", X"00000000000000000000000000000000", X"EDC58173B381AC54D86D7334E069924F"),
    (X"F8000000000000000000000000000000", X"00000000000000000000000000000000", X"2AE2B1FBF8DAE9D3F2E9ECF96B8EA287"),
    (X"FC000000000000000000000000000000", X"00000000000000000000000000000000", X"855A70CBCA780A83D4AEDE10206FD117"),
    (X"FE000000000000000000000000000000", X"00000000000000000000000000000000", X"1A625E640BDC50FB10936C1C1C3FBE88"),
    (X"FF000000000000000000000000000000", X"00000000000000000000000000000000", X"83EA834DED44FDF795DF4B189B5EB8F5"),
    (X"FF800000000000000000000000000000", X"00000000000000000000000000000000", X"D88D500984FE9A8DA0BF891DA2AB67D1"),
    (X"FFC00000000000000000000000000000", X"00000000000000000000000000000000", X"44B43BB05F1DFAE3682448FF9B809BDE"),
    (X"FFE00000000000000000000000000000", X"00000000000000000000000000000000", X"C2DB48B274F0BA91BB5E5EC624FBEC06"),
    (X"FFF00000000000000000000000000000", X"00000000000000000000000000000000", X"E575E7B0C46AEE8C19902C075406C358"),
    (X"FFF80000000000000000000000000000", X"00000000000000000000000000000000", X"FC04B70C143A3FF003B05EADFA1FC24A"),
    (X"FFFC0000000000000000000000000000", X"00000000000000000000000000000000", X"B8FA48ADC05916A36A739A3C639CC5F9"),
    (X"FFFE0000000000000000000000000000", X"00000000000000000000000000000000", X"14A50D987D23278977F1266AC2DC5F6C"),
    (X"FFFF0000000000000000000000000000", X"00000000000000000000000000000000", X"62980269B1A94C6C97B3A53720B440A2"),
    (X"FFFF8000000000000000000000000000", X"00000000000000000000000000000000", X"400B76B5778D1842CBE3329B63B9DE74"),
    (X"FFFFC000000000000000000000000000", X"00000000000000000000000000000000", X"430AE287C864D59EC66BF78D95FB0169"),
    (X"FFFFE000000000000000000000000000", X"00000000000000000000000000000000", X"E5F30592466A8C89611B028688C451AC"),
    (X"FFFFF000000000000000000000000000", X"00000000000000000000000000000000", X"A830081AD40DAB53DBAFD4B4A0A976A8"),
    (X"FFFFF800000000000000000000000000", X"00000000000000000000000000000000", X"F5713B8D952DCA4CC023B3C3230963BA"),
    (X"FFFFFC00000000000000000000000000", X"00000000000000000000000000000000", X"90DC21D7B4E9AA0E9F4789AD10BCC779"),
    (X"FFFFFE00000000000000000000000000", X"00000000000000000000000000000000", X"BFF8E0F1F2ADBBA39EBBFC833FAF41F9"),
    (X"FFFFFF00000000000000000000000000", X"00000000000000000000000000000000", X"C016046DD57AA2D9937846F5BDCBC222"),
    (X"FFFFFF80000000000000000000000000", X"00000000000000000000000000000000", X"0442DDAE7D6776DE59F12804D16EE82F"),
    (X"FFFFFFC0000000000000000000000000", X"00000000000000000000000000000000", X"BD878C6D00CCDAEE21EE6A67AC67363E"),
    (X"FFFFFFE0000000000000000000000000", X"00000000000000000000000000000000", X"777EA3A77C12022F8976299C8ED7774A"),
    (X"FFFFFFF0000000000000000000000000", X"00000000000000000000000000000000", X"E5DCF13452D899C0F9B18DB44A0F3A5A"),
    (X"FFFFFFF8000000000000000000000000", X"00000000000000000000000000000000", X"9C3B4689A65081F6D98E30EDE67B08E9"),
    (X"FFFFFFFC000000000000000000000000", X"00000000000000000000000000000000", X"48D36CBB7C7C110CAE598DDD5C9B4999"),
    (X"FFFFFFFE000000000000000000000000", X"00000000000000000000000000000000", X"44D34C4A4C9133ABB3E31D7B33BCE5CF"),
    (X"FFFFFFFF000000000000000000000000", X"00000000000000000000000000000000", X"E910C7E0E49DA858B58404A9B4331C95"),
    (X"FFFFFFFF800000000000000000000000", X"00000000000000000000000000000000", X"4026B5DFED768FEBF2D4934D66B8F91E"),
    (X"FFFFFFFFC00000000000000000000000", X"00000000000000000000000000000000", X"E12F718CF6E289DDB3B6D743DC833F2F"),
    (X"FFFFFFFFE00000000000000000000000", X"00000000000000000000000000000000", X"6F81DACA6CF40DDA1310582377FC68D8"),
    (X"FFFFFFFFF00000000000000000000000", X"00000000000000000000000000000000", X"35E568A20A49B3739DF495F42AB6389B"),
    (X"FFFFFFFFF80000000000000000000000", X"00000000000000000000000000000000", X"AF1019A2448F186124AA1A4C43B9D803"),
    (X"FFFFFFFFFC0000000000000000000000", X"00000000000000000000000000000000", X"57162D1025A79438001F60C82727C9E9"),
    (X"FFFFFFFFFE0000000000000000000000", X"00000000000000000000000000000000", X"1F6E7D6CB5F9EDDFB4DD407ABFAF5C89"),
    (X"FFFFFFFFFF0000000000000000000000", X"00000000000000000000000000000000", X"D92F1CC823A93FAC4540303CA9F93269"),
    (X"FFFFFFFFFF8000000000000000000000", X"00000000000000000000000000000000", X"9183BD80A1F6FC759AB3428E5D7D0A9C"),
    (X"FFFFFFFFFFC000000000000000000000", X"00000000000000000000000000000000", X"37610DD9EC7AD6371A05A87364371144"),
    (X"FFFFFFFFFFE000000000000000000000", X"00000000000000000000000000000000", X"827D0941F270ACED90BB4CDD7B8E24C0"),
    (X"FFFFFFFFFFF000000000000000000000", X"00000000000000000000000000000000", X"A60C67A52E34F585C35A149354F65A6D"),
    (X"FFFFFFFFFFF800000000000000000000", X"00000000000000000000000000000000", X"EF9343F30261DF3AB616F6B6F08E3E94"),
    (X"FFFFFFFFFFFC00000000000000000000", X"00000000000000000000000000000000", X"D3EA7C59822CD6AD5DFD1D74059BF50C"),
    (X"FFFFFFFFFFFE00000000000000000000", X"00000000000000000000000000000000", X"2BA6F2E165099874D4908E96F85CFA9C"),
    (X"FFFFFFFFFFFF00000000000000000000", X"00000000000000000000000000000000", X"7F751EF0100DDFC081630872A23B4607"),
    (X"FFFFFFFFFFFF80000000000000000000", X"00000000000000000000000000000000", X"B899D9BF6F6BFFEBF1F4FDCC5C631E20"),
    (X"FFFFFFFFFFFFC0000000000000000000", X"00000000000000000000000000000000", X"ECEBB8D8F8952A9EB79E649A7E7802FA"),
    (X"FFFFFFFFFFFFE0000000000000000000", X"00000000000000000000000000000000", X"ACAE850E3ECDE60A1B59B31C88613740"),
    (X"FFFFFFFFFFFFF0000000000000000000", X"00000000000000000000000000000000", X"F2D6128327C86833987EC81F9F9F6E34"),
    (X"FFFFFFFFFFFFF8000000000000000000", X"00000000000000000000000000000000", X"F537D7E25603BA4A52EE65345014122D"),
    (X"FFFFFFFFFFFFFC000000000000000000", X"00000000000000000000000000000000", X"E10D7D4A9C678BAD6B5888F6E9765231"),
    (X"FFFFFFFFFFFFFE000000000000000000", X"00000000000000000000000000000000", X"02494307793210504C75A06080672F71"),
    (X"FFFFFFFFFFFFFF000000000000000000", X"00000000000000000000000000000000", X"A0A95F87B535416335A5C232971AF785"),
    (X"FFFFFFFFFFFFFF800000000000000000", X"00000000000000000000000000000000", X"1E627F8148E5B068DF50DEA0DD6218EB"),
    (X"FFFFFFFFFFFFFFC00000000000000000", X"00000000000000000000000000000000", X"60198C0F74EE1E2AA3B1415401A45FC1"),
    (X"FFFFFFFFFFFFFFE00000000000000000", X"00000000000000000000000000000000", X"1526964A1CB7AB50E03EEE638AA3C0EA"),
    (X"FFFFFFFFFFFFFFF00000000000000000", X"00000000000000000000000000000000", X"10A5A84D3929AC60114089718EFFE7A5"),
    (X"FFFFFFFFFFFFFFF80000000000000000", X"00000000000000000000000000000000", X"7AB8F889D71E00F9A35E005DADA154F6"),
    (X"FFFFFFFFFFFFFFFC0000000000000000", X"00000000000000000000000000000000", X"7DB29053292918072667700F1568DDF9"),
    (X"FFFFFFFFFFFFFFFE0000000000000000", X"00000000000000000000000000000000", X"975FA30DB8808D2D0B55A63D77886440"),
    (X"FFFFFFFFFFFFFFFF0000000000000000", X"00000000000000000000000000000000", X"F9479211DA0BD50FAEE83F1565830BB8"),
    (X"FFFFFFFFFFFFFFFF8000000000000000", X"00000000000000000000000000000000", X"9F1F6B5762EA741952F9E780833C281C"),
    (X"FFFFFFFFFFFFFFFFC000000000000000", X"00000000000000000000000000000000", X"C48F3A601C22448E6F52A0C6C58CC6A3"),
    (X"FFFFFFFFFFFFFFFFE000000000000000", X"00000000000000000000000000000000", X"5111EA5FDDB6A22F2C7D6A501372EC05"),
    (X"FFFFFFFFFFFFFFFFF000000000000000", X"00000000000000000000000000000000", X"0D39C870F3D7C25698449BC3A523978A"),
    (X"FFFFFFFFFFFFFFFFF800000000000000", X"00000000000000000000000000000000", X"B9636FECA0D3D73D7376D27ADDF3A6AC"),
    (X"FFFFFFFFFFFFFFFFFC00000000000000", X"00000000000000000000000000000000", X"79C61AE1E6BFF595752EFC86100524DD"),
    (X"FFFFFFFFFFFFFFFFFE00000000000000", X"00000000000000000000000000000000", X"F95518B35556EB3462FE23350287B32C"),
    (X"FFFFFFFFFFFFFFFFFF00000000000000", X"00000000000000000000000000000000", X"CF8F7F8920C804914F2234B60BBD9DA5"),
    (X"FFFFFFFFFFFFFFFFFF80000000000000", X"00000000000000000000000000000000", X"4FB50BC022141EE6838E8C9185D52076"),
    (X"FFFFFFFFFFFFFFFFFFC0000000000000", X"00000000000000000000000000000000", X"92EBBDC0E8EBE02D8D6C0B70263D503A"),
    (X"FFFFFFFFFFFFFFFFFFE0000000000000", X"00000000000000000000000000000000", X"9C5D80FAEB4CB0B6773E428C2BDF0110"),
    (X"FFFFFFFFFFFFFFFFFFF0000000000000", X"00000000000000000000000000000000", X"90E61074CDE1BAAF424AD2301E0058CA"),
    (X"FFFFFFFFFFFFFFFFFFF8000000000000", X"00000000000000000000000000000000", X"8C3078D7FAF6F1B51D9097EE86F96BDD"),
    (X"FFFFFFFFFFFFFFFFFFFC000000000000", X"00000000000000000000000000000000", X"E9CD8772692C5C6A8295F32E786D8F3A"),
    (X"FFFFFFFFFFFFFFFFFFFE000000000000", X"00000000000000000000000000000000", X"1C2732B3DCD061EFA2E3FFA4BD84CA47"),
    (X"FFFFFFFFFFFFFFFFFFFF000000000000", X"00000000000000000000000000000000", X"FADE2B6970BDE3F443FEF947208D9FFF"),
    (X"FFFFFFFFFFFFFFFFFFFF800000000000", X"00000000000000000000000000000000", X"A526F811EDA6553BD45FC862AFC1AA05"),
    (X"FFFFFFFFFFFFFFFFFFFFC00000000000", X"00000000000000000000000000000000", X"7FE38E8821D1CCA02DFC7F3B090CF0ED"),
    (X"FFFFFFFFFFFFFFFFFFFFE00000000000", X"00000000000000000000000000000000", X"678D8AA0257AE752A69D5FC231CDBFB5"),
    (X"FFFFFFFFFFFFFFFFFFFFF00000000000", X"00000000000000000000000000000000", X"3F015B261B4729C211035507729D0578"),
    (X"FFFFFFFFFFFFFFFFFFFFF80000000000", X"00000000000000000000000000000000", X"D7C894C022FC515F14164F6BB1BB7B00"),
    (X"FFFFFFFFFFFFFFFFFFFFFC0000000000", X"00000000000000000000000000000000", X"3F7D7274917CCEB3EFFA7247238A9444"),
    (X"FFFFFFFFFFFFFFFFFFFFFE0000000000", X"00000000000000000000000000000000", X"02795B3F04DBA054A73C57CBACDB284B"),
    (X"FFFFFFFFFFFFFFFFFFFFFF0000000000", X"00000000000000000000000000000000", X"4A7934672C16654C7544D92050CB9F3D"),
    (X"FFFFFFFFFFFFFFFFFFFFFF8000000000", X"00000000000000000000000000000000", X"012F2E4D901CE0B96DA7F0CDB2908259"),
    (X"FFFFFFFFFFFFFFFFFFFFFFC000000000", X"00000000000000000000000000000000", X"D9C34EE50CF33FDDB9102CFA8DAF4322"),
    (X"FFFFFFFFFFFFFFFFFFFFFFE000000000", X"00000000000000000000000000000000", X"E39BA037293D377BB16A4699917D1F70"),
    (X"FFFFFFFFFFFFFFFFFFFFFFF000000000", X"00000000000000000000000000000000", X"05C3890964B37EE2DE7984A7CDC5A968"),
    (X"FFFFFFFFFFFFFFFFFFFFFFF800000000", X"00000000000000000000000000000000", X"AA32D893D73A538571C4E1ECA0496467"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFC00000000", X"00000000000000000000000000000000", X"99DBDBF5A773921BAC712690688CF676"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFE00000000", X"00000000000000000000000000000000", X"EC482A5705E45A05770F19C943EC37B2"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFF00000000", X"00000000000000000000000000000000", X"CC64CD1C2CBAA529446DA6406C94EC51"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFF80000000", X"00000000000000000000000000000000", X"E8A86E3D2A3FC225D8033749AACA3BF2"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000", X"00000000000000000000000000000000", X"406B87BA4AA0F141039DBE915A2B3348"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000", X"00000000000000000000000000000000", X"935B7103DEF16EB8D8B79CFD0DC1A134"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000", X"00000000000000000000000000000000", X"B5529D9BE0131D8215DD65C4E34630A2"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000", X"00000000000000000000000000000000", X"933B62A5760672686B3D6062B6180D6B"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000", X"00000000000000000000000000000000", X"940A9886821A5B0E7D15BEEA65F242A6"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000", X"00000000000000000000000000000000", X"D372A141E86D3F3224D6150860ABD01A"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000", X"00000000000000000000000000000000", X"8AD229B568F51B744F7842B1FE9AE188"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000", X"00000000000000000000000000000000", X"6B4E294FFAED07E7278E539A1A6985C9"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000", X"00000000000000000000000000000000", X"B2E9D35B0AD46CF1ACEECFE49FE8527A"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000", X"00000000000000000000000000000000", X"5C40CF411B315751B2A032334D2E9417"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000", X"00000000000000000000000000000000", X"B80B9D8094340CAE0E2FE4525A847222"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000", X"00000000000000000000000000000000", X"E4C07D628EB21E39F2BA1B5340A18E13"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000", X"00000000000000000000000000000000", X"835A1E7D79A283F02E082FEF5946EAA1"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000", X"00000000000000000000000000000000", X"7AD2E9FBA2B913B763405D44D520643D"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000", X"00000000000000000000000000000000", X"E5D224A228BBD5BE80C255BB63AD854A"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000", X"00000000000000000000000000000000", X"493CC65C8C65EE3EC2E7FEB1F2E2688D"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000", X"00000000000000000000000000000000", X"A36C6BDA232148E0844189B34A0645E0"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000", X"00000000000000000000000000000000", X"4E3A57CFDCC9C9DA0D774F073029DB28"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000", X"00000000000000000000000000000000", X"C9D5B2EE3292B262A79192BB81107006"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800", X"00000000000000000000000000000000", X"A1DDB1C43BC3DF36F0A23FE88E9A7DCA"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00", X"00000000000000000000000000000000", X"D237DB2C37BBC6189ADEC6E4612B38F5"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00", X"00000000000000000000000000000000", X"EA459A91531D5B98211C81B43644E370"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00", X"00000000000000000000000000000000", X"EB6B8A389564056730B7569C0C855D3E"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80", X"00000000000000000000000000000000", X"77C6322B360ACFFB464FD8A5AED6AA47"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0", X"00000000000000000000000000000000", X"8ED8E0FC0E95A6746385F52F7D8DCB4E"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0", X"00000000000000000000000000000000", X"E15A4D5D1D47B8231D4ADD95FECFAB70"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0", X"00000000000000000000000000000000", X"F3A87234260FFDAFD9065555AA0CDABA"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8", X"00000000000000000000000000000000", X"32BB535356C6519479AECCD8328DD064"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC", X"00000000000000000000000000000000", X"EF49C8F00D3DBD7340A7F55784A81BB8"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE", X"00000000000000000000000000000000", X"6423F8EF0E060342865611718B62D49B"),
    (X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF", X"00000000000000000000000000000000", X"952ABAC4EBDA6CE9D1CAE8F2639F2B74")
    );
end package aesTest_GRBC_s18;
