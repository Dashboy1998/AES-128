use work.data_types.all;

package rcon_table is
	constant rcon_LUT : AByte := (X"B1",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"1B",X"36");
end rcon_table;