use work.data_types.all;

entity multVector is
	port(
	A: in word;
	