use work.LUT_array.all;

package LUT2_array is
	type array_512 is array (0 to 1) of array_256;
end LUT2_array;