library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package aes128Test is
  type test is record
    key      : std_logic_vector(0 to 127);
    plain    : std_logic_vector(0 to 127);
    expected : std_logic_vector(0 to 127);
  end record test;
  type testArray is array (natural range <>) of test;
  constant tests : testarray := (
	(X"000102030405060708090A0B0C0D0E0F", X"00112233445566778899AABBCCDDEEFF", X"69C4E0D86A7B0430D8CDB78070B4C55A"),
    (X"00000000000000000000000000000000", X"80000000000000000000000000000000", X"3AD78E726C1EC02B7EBFE92B23D9EC34"),
	(X"00000000000000000000000000000000", X"C0000000000000000000000000000000", X"AAE5939C8EFDF2F04E60B9FE7117B2C2"),
	(X"00000000000000000000000000000000", X"E0000000000000000000000000000000", X"F031D4D74F5DCBF39DAAF8CA3AF6E527"),
	(X"00000000000000000000000000000000", X"F0000000000000000000000000000000", X"96D9FD5CC4F07441727DF0F33E401A36"),
	(X"00000000000000000000000000000000", X"F8000000000000000000000000000000", X"30CCDB044646D7E1F3CCEA3DCA08B8C0"),
	(X"00000000000000000000000000000000", X"FC000000000000000000000000000000", X"16AE4CE5042A67EE8E177B7C587ECC82"),
	(X"00000000000000000000000000000000", X"FE000000000000000000000000000000", X"B6DA0BB11A23855D9C5CB1B4C6412E0A"),
	(X"00000000000000000000000000000000", X"FF000000000000000000000000000000", X"DB4F1AA530967D6732CE4715EB0EE24B"),
	(X"00000000000000000000000000000000", X"FF800000000000000000000000000000", X"A81738252621DD180A34F3455B4BAA2F"),
	(X"00000000000000000000000000000000", X"FFC00000000000000000000000000000", X"77E2B508DB7FD89234CAF7939EE5621A"),
	(X"00000000000000000000000000000000", X"FFE00000000000000000000000000000", X"B8499C251F8442EE13F0933B688FCD19"),
	(X"00000000000000000000000000000000", X"FFF00000000000000000000000000000", X"965135F8A81F25C9D630B17502F68E53"),
	(X"00000000000000000000000000000000", X"FFF80000000000000000000000000000", X"8B87145A01AD1C6CEDE995EA3670454F"),
	(X"00000000000000000000000000000000", X"FFFC0000000000000000000000000000", X"8EAE3B10A0C8CA6D1D3B0FA61E56B0B2"),
	(X"00000000000000000000000000000000", X"FFFE0000000000000000000000000000", X"64B4D629810FDA6BAFDF08F3B0D8D2C5"),
	(X"00000000000000000000000000000000", X"FFFF0000000000000000000000000000", X"D7E5DBD3324595F8FDC7D7C571DA6C2A"),
	(X"00000000000000000000000000000000", X"FFFF8000000000000000000000000000", X"F3F72375264E167FCA9DE2C1527D9606"),
	(X"00000000000000000000000000000000", X"FFFFC000000000000000000000000000", X"8EE79DD4F401FF9B7EA945D86666C13B"),
	(X"00000000000000000000000000000000", X"FFFFE000000000000000000000000000", X"DD35CEA2799940B40DB3F819CB94C08B"),
	(X"00000000000000000000000000000000", X"FFFFF000000000000000000000000000", X"6941CB6B3E08C2B7AFA581EBDD607B87"),
	(X"00000000000000000000000000000000", X"FFFFF800000000000000000000000000", X"2C20F439F6BB097B29B8BD6D99AAD799"),
	(X"00000000000000000000000000000000", X"FFFFFC00000000000000000000000000", X"625D01F058E565F77AE86378BD2C49B3"),
	(X"00000000000000000000000000000000", X"FFFFFE00000000000000000000000000", X"C0B5FD98190EF45FBB4301438D095950"),
	(X"00000000000000000000000000000000", X"FFFFFF00000000000000000000000000", X"13001FF5D99806EFD25DA34F56BE854B"),
	(X"00000000000000000000000000000000", X"FFFFFF80000000000000000000000000", X"3B594C60F5C8277A5113677F94208D82"),
	(X"00000000000000000000000000000000", X"FFFFFFC0000000000000000000000000", X"E9C0FC1818E4AA46BD2E39D638F89E05"),
	(X"00000000000000000000000000000000", X"FFFFFFE0000000000000000000000000", X"F8023EE9C3FDC45A019B4E985C7E1A54"),
	(X"00000000000000000000000000000000", X"FFFFFFF0000000000000000000000000", X"35F40182AB4662F3023BAEC1EE796B57"),
	(X"00000000000000000000000000000000", X"FFFFFFF8000000000000000000000000", X"3AEBBAD7303649B4194A6945C6CC3694"),
	(X"00000000000000000000000000000000", X"FFFFFFFC000000000000000000000000", X"A2124BEA53EC2834279BED7F7EB0F938"),
	(X"00000000000000000000000000000000", X"FFFFFFFE000000000000000000000000", X"B9FB4399FA4FACC7309E14EC98360B0A"),
	(X"00000000000000000000000000000000", X"FFFFFFFF000000000000000000000000", X"C26277437420C5D634F715AEA81A9132"),
	(X"00000000000000000000000000000000", X"FFFFFFFF800000000000000000000000", X"171A0E1B2DD424F0E089AF2C4C10F32F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFC00000000000000000000000", X"7CADBE402D1B208FE735EDCE00AEE7CE"),
	(X"00000000000000000000000000000000", X"FFFFFFFFE00000000000000000000000", X"43B02FF929A1485AF6F5C6D6558BAA0F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFF00000000000000000000000", X"092FAACC9BF43508BF8FA8613CA75DEA"),
	(X"00000000000000000000000000000000", X"FFFFFFFFF80000000000000000000000", X"CB2BF8280F3F9742C7ED513FE802629C"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFC0000000000000000000000", X"215A41EE442FA992A6E323986DED3F68"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFE0000000000000000000000", X"F21E99CF4F0F77CEA836E11A2FE75FB1"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFF0000000000000000000000", X"95E3A0CA9079E646331DF8B4E70D2CD6"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFF8000000000000000000000", X"4AFE7F120CE7613F74FC12A01A828073"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFC000000000000000000000", X"827F000E75E2C8B9D479BEED913FE678"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFE000000000000000000000", X"35830C8E7AAEFE2D30310EF381CBF691"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFF000000000000000000000", X"191AA0F2C8570144F38657EA4085EBE5"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFF800000000000000000000", X"85062C2C909F15D9269B6C18CE99C4F0"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFC00000000000000000000", X"678034DC9E41B5A560ED239EEAB1BC78"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFE00000000000000000000", X"C2F93A4CE5AB6D5D56F1B93CF19911C1"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFF00000000000000000000", X"1C3112BCB0C1DCC749D799743691BF82"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFF80000000000000000000", X"00C55BD75C7F9C881989D3EC1911C0D4"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFC0000000000000000000", X"EA2E6B5EF182B7DFF3629ABD6A12045F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFE0000000000000000000", X"22322327E01780B17397F24087F8CC6F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFF0000000000000000000", X"C9CACB5CD11692C373B2411768149EE7"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFF8000000000000000000", X"A18E3DBBCA577860DAB6B80DA3139256"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFC000000000000000000", X"79B61C37BF328ECCA8D743265A3D425C"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFE000000000000000000", X"D2D99C6BCC1F06FDA8E27E8AE3F1CCC7"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFF000000000000000000", X"1BFD4B91C701FD6B61B7F997829D663B"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFF800000000000000000", X"11005D52F25F16BDC9545A876A63490A"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFC00000000000000000", X"3A4D354F02BB5A5E47D39666867F246A"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFE00000000000000000", X"D451B8D6E1E1A0EBB155FBBF6E7B7DC3"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFF00000000000000000", X"6898D4F42FA7BA6A10AC05E87B9F2080"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFF80000000000000000", X"B611295E739CA7D9B50F8E4C0E754A3F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFC0000000000000000", X"7D33FC7D8ABE3CA1936759F8F5DEAF20"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFE0000000000000000", X"3B5E0F566DC96C298F0C12637539B25C"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFF0000000000000000", X"F807C3E7985FE0F5A50E2CDB25C5109E"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFF8000000000000000", X"41F992A856FB278B389A62F5D274D7E9"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFC000000000000000", X"10D3ED7A6FE15AB4D91ACBC7D0767AB1"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFE000000000000000", X"21FEECD45B2E675973AC33BF0C5424FC"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFF000000000000000", X"1480CB3955BA62D09EEA668F7C708817"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFF800000000000000", X"66404033D6B72B609354D5496E7EB511"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFC00000000000000", X"1C317A220A7D700DA2B1E075B00266E1"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFE00000000000000", X"AB3B89542233F1271BF8FD0C0F403545"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFF00000000000000", X"D93EAE966FAC46DCA927D6B114FA3F9E"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFF80000000000000", X"1BDEC521316503D9D5EE65DF3EA94DDF"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFC0000000000000", X"EEF456431DEA8B4ACF83BDAE3717F75F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFE0000000000000", X"06F2519A2FAFAA596BFEF5CFA15C21B9"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFF0000000000000", X"251A7EAC7E2FE809E4AA8D0D7012531A"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFF8000000000000", X"3BFFC16E4C49B268A20F8D96A60B4058"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFC000000000000", X"E886F9281999C5BB3B3E8862E2F7C988"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFE000000000000", X"563BF90D61BEEF39F48DD625FCEF1361"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFF000000000000", X"4D37C850644563C69FD0ACD9A049325B"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFF800000000000", X"B87C921B91829EF3B13CA541EE1130A6"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFC00000000000", X"2E65EB6B6EA383E109ACCCE8326B0393"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFE00000000000", X"9CA547F7439EDC3E255C0F4D49AA8990"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFF00000000000", X"A5E652614C9300F37816B1F9FD0C87F9"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFF80000000000", X"14954F0B4697776F44494FE458D814ED"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFC0000000000", X"7C8D9AB6C2761723FE42F8BB506CBCF7"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFE0000000000", X"DB7E1932679FDD99742AAB04AA0D5A80"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFF0000000000", X"4C6A1C83E568CD10F27C2D73DED19C28"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFF8000000000", X"90ECBE6177E674C98DE412413F7AC915"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFC000000000", X"90684A2AC55FE1EC2B8EBD5622520B73"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFE000000000", X"7472F9A7988607CA79707795991035E6"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFF000000000", X"56AFF089878BF3352F8DF172A3AE47D8"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFF800000000", X"65C0526CBE40161B8019A2A3171ABD23"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFC00000000", X"377BE0BE33B4E3E310B4AABDA173F84F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFE00000000", X"9402E9AA6F69DE6504DA8D20C4FCAA2F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFF00000000", X"123C1F4AF313AD8C2CE648B2E71FB6E1"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFF80000000", X"1FFC626D30203DCDB0019FB80F726CF4"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000", X"76DA1FBE3A50728C50FD2E621B5AD885"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000", X"082EB8BE35F442FB52668E16A591D1D6"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000", X"E656F9ECF5FE27EC3E4A73D00C282FB3"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000", X"2CA8209D63274CD9A29BB74BCD77683A"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000", X"79BF5DCE14BB7DD73A8E3611DE7CE026"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000", X"3C849939A5D29399F344C4A0ECA8A576"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000", X"ED3C0A94D59BECE98835DA7AA4F07CA2"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000", X"63919ED4CE10196438B6AD09D99CD795"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000", X"7678F3A833F19FEA95F3C6029E2BC610"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000", X"3AA426831067D36B92BE7C5F81C13C56"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000", X"9272E2D2CDD11050998C845077A30EA0"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000", X"088C4B53F5EC0FF814C19ADAE7F6246C"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000", X"4010A5E401FDF0A0354DDBCC0D012B17"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000", X"A87A385736C0A6189BD6589BD8445A93"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000", X"545F2B83D9616DCCF60FA9830E9CD287"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000", X"4B706F7F92406352394037A6D4F4688D"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000", X"B7972B3941C44B90AFA7B264BFBA7387"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000", X"6F45732CF10881546F0FD23896D2BB60"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000", X"2E3579CA15AF27F64B3C955A5BFC30BA"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800", X"34A2C5A91AE2AEC99B7D1B5FA6780447"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00", X"A4D6616BD04F87335B0E53351227A9EE"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00", X"7F692B03945867D16179A8CEFC83EA3F"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00", X"3BD141EE84A0E6414A26E7A4F281F8A2"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80", X"D1788F572D98B2B16EC5D5F3922B99BC"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0", X"0833FF6F61D98A57B288E8C3586B85A6"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0", X"8568261797DE176BF0B43BECC6285AFB"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0", X"F9B0FDA0C4A898F5B9E6F661C4CE4D07"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8", X"8ADE895913685C67C5269F8AAE42983E"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC", X"39BDE67D5C8ED8A8B1C37EB8FA9F5AC0"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE", X"5C005E72C1418C44F569F2EA33BA54F3"),
	(X"00000000000000000000000000000000", X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF", X"3F5B8CC9EA855A0AFA7347D23E8D664E"),
	(X"80000000000000000000000000000000", X"00000000000000000000000000000000", X"0EDD33D3C621E546455BD8BA1418BEC8"),
	(X"C0000000000000000000000000000000", X"00000000000000000000000000000000", X"4BC3F883450C113C64CA42E1112A9E87"),
	(X"E0000000000000000000000000000000", X"00000000000000000000000000000000", X"72A1DA770F5D7AC4C9EF94D822AFFD97"),
	(X"F0000000000000000000000000000000", X"00000000000000000000000000000000", X"970014D634E2B7650777E8E84D03CCD8"),
	(X"F8000000000000000000000000000000", X"00000000000000000000000000000000", X"F17E79AED0DB7E279E955B5F493875A7"),
	(X"FC000000000000000000000000000000", X"00000000000000000000000000000000", X"9ED5A75136A940D0963DA379DB4AF26A"),
	(X"FE000000000000000000000000000000", X"00000000000000000000000000000000", X"C4295F83465C7755E8FA364BAC6A7EA5"),
	(X"FF000000000000000000000000000000", X"00000000000000000000000000000000", X"B1D758256B28FD850AD4944208CF1155"),
	(X"FF800000000000000000000000000000", X"00000000000000000000000000000000", X"42FFB34C743DE4D88CA38011C990890B"),
	(X"FFC00000000000000000000000000000", X"00000000000000000000000000000000", X"9958F0ECEA8B2172C0C1995F9182C0F3"),
	(X"FFE00000000000000000000000000000", X"00000000000000000000000000000000", X"956D7798FAC20F82A8823F984D06F7F5"),
	(X"FFF00000000000000000000000000000", X"00000000000000000000000000000000", X"A01BF44F2D16BE928CA44AAF7B9B106B"),
	(X"FFF80000000000000000000000000000", X"00000000000000000000000000000000", X"B5F1A33E50D40D103764C76BD4C6B6F8"),
	(X"FFFC0000000000000000000000000000", X"00000000000000000000000000000000", X"2637050C9FC0D4817E2D69DE878AEE8D"),
	(X"FFFE0000000000000000000000000000", X"00000000000000000000000000000000", X"113ECBE4A453269A0DD26069467FB5B5"),
	(X"FFFF0000000000000000000000000000", X"00000000000000000000000000000000", X"97D0754FE68F11B9E375D070A608C884"),
	(X"FFFF8000000000000000000000000000", X"00000000000000000000000000000000", X"C6A0B3E998D05068A5399778405200B4"),
	(X"FFFFC000000000000000000000000000", X"00000000000000000000000000000000", X"DF556A33438DB87BC41B1752C55E5E49"),
	(X"FFFFE000000000000000000000000000", X"00000000000000000000000000000000", X"90FB128D3A1AF6E548521BB962BF1F05"),
	(X"FFFFF000000000000000000000000000", X"00000000000000000000000000000000", X"26298E9C1DB517C215FADFB7D2A8D691"),
	(X"FFFFF800000000000000000000000000", X"00000000000000000000000000000000", X"A6CB761D61F8292D0DF393A279AD0380"),
	(X"FFFFFC00000000000000000000000000", X"00000000000000000000000000000000", X"12ACD89B13CD5F8726E34D44FD486108"),
	(X"FFFFFE00000000000000000000000000", X"00000000000000000000000000000000", X"95B1703FC57BA09FE0C3580FEBDD7ED4"),
	(X"FFFFFF00000000000000000000000000", X"00000000000000000000000000000000", X"DE11722D893E9F9121C381BECC1DA59A"),
	(X"FFFFFF80000000000000000000000000", X"00000000000000000000000000000000", X"6D114CCB27BF391012E8974C546D9BF2"),
	(X"FFFFFFC0000000000000000000000000", X"00000000000000000000000000000000", X"5CE37E17EB4646ECFAC29B9CC38D9340"),
	(X"FFFFFFE0000000000000000000000000", X"00000000000000000000000000000000", X"18C1B6E2157122056D0243D8A165CDDB"),
	(X"FFFFFFF0000000000000000000000000", X"00000000000000000000000000000000", X"99693E6A59D1366C74D823562D7E1431"),
	(X"FFFFFFF8000000000000000000000000", X"00000000000000000000000000000000", X"6C7C64DC84A8BBA758ED17EB025A57E3"),
	(X"FFFFFFFC000000000000000000000000", X"00000000000000000000000000000000", X"E17BC79F30EAAB2FAC2CBBE3458D687A"),
	(X"FFFFFFFE000000000000000000000000", X"00000000000000000000000000000000", X"1114BC2028009B923F0B01915CE5E7C4"),
	(X"FFFFFFFF000000000000000000000000", X"00000000000000000000000000000000", X"9C28524A16A1E1C1452971CAA8D13476"),
	(X"FFFFFFFF800000000000000000000000", X"00000000000000000000000000000000", X"ED62E16363638360FDD6AD62112794F0"),
	(X"FFFFFFFFC00000000000000000000000", X"00000000000000000000000000000000", X"5A8688F0B2A2C16224C161658FFD4044"),
	(X"FFFFFFFFE00000000000000000000000", X"00000000000000000000000000000000", X"23F710842B9BB9C32F26648C786807CA"),
	(X"FFFFFFFFF00000000000000000000000", X"00000000000000000000000000000000", X"44A98BF11E163F632C47EC6A49683A89"),
	(X"FFFFFFFFF80000000000000000000000", X"00000000000000000000000000000000", X"0F18AFF94274696D9B61848BD50AC5E5"),
	(X"FFFFFFFFFC0000000000000000000000", X"00000000000000000000000000000000", X"82408571C3E2424540207F833B6DDA69"),
	(X"FFFFFFFFFE0000000000000000000000", X"00000000000000000000000000000000", X"303FF996947F0C7D1F43C8F3027B9B75"),
	(X"FFFFFFFFFF0000000000000000000000", X"00000000000000000000000000000000", X"7DF4DAF4AD29A3615A9B6ECE5C99518A"),
	(X"FFFFFFFFFF8000000000000000000000", X"00000000000000000000000000000000", X"C72954A48D0774DB0B4971C526260415"),
	(X"FFFFFFFFFFC000000000000000000000", X"00000000000000000000000000000000", X"1DF9B76112DC6531E07D2CFDA04411F0"),
	(X"FFFFFFFFFFE000000000000000000000", X"00000000000000000000000000000000", X"8E4D8E699119E1FC87545A647FB1D34F"),
	(X"FFFFFFFFFFF000000000000000000000", X"00000000000000000000000000000000", X"E6C4807AE11F36F091C57D9FB68548D1"),
	(X"FFFFFFFFFFF800000000000000000000", X"00000000000000000000000000000000", X"8EBF73AAD49C82007F77A5C1CCEC6AB4"),
	(X"FFFFFFFFFFFC00000000000000000000", X"00000000000000000000000000000000", X"4FB288CC2040049001D2C7585AD123FC"),
	(X"FFFFFFFFFFFE00000000000000000000", X"00000000000000000000000000000000", X"04497110EFB9DCEB13E2B13FB4465564"),
	(X"FFFFFFFFFFFF00000000000000000000", X"00000000000000000000000000000000", X"75550E6CB5A88E49634C9AB69EDA0430"),
	(X"FFFFFFFFFFFF80000000000000000000", X"00000000000000000000000000000000", X"B6768473CE9843EA66A81405DD50B345"),
	(X"FFFFFFFFFFFFC0000000000000000000", X"00000000000000000000000000000000", X"CB2F430383F9084E03A653571E065DE6"),
	(X"FFFFFFFFFFFFE0000000000000000000", X"00000000000000000000000000000000", X"FF4E66C07BAE3E79FB7D210847A3B0BA"),
	(X"FFFFFFFFFFFFF0000000000000000000", X"00000000000000000000000000000000", X"7B90785125505FAD59B13C186DD66CE3"),
	(X"FFFFFFFFFFFFF8000000000000000000", X"00000000000000000000000000000000", X"8B527A6AEBDAEC9EAEF8EDA2CB7783E5"),
	(X"FFFFFFFFFFFFFC000000000000000000", X"00000000000000000000000000000000", X"43FDAF53EBBC9880C228617D6A9B548B"),
	(X"FFFFFFFFFFFFFE000000000000000000", X"00000000000000000000000000000000", X"53786104B9744B98F052C46F1C850D0B"),
	(X"FFFFFFFFFFFFFF000000000000000000", X"00000000000000000000000000000000", X"B5AB3013DD1E61DF06CBAF34CA2AEE78"),
	(X"FFFFFFFFFFFFFF800000000000000000", X"00000000000000000000000000000000", X"7470469BE9723030FDCC73A8CD4FBB10"),
	(X"FFFFFFFFFFFFFFC00000000000000000", X"00000000000000000000000000000000", X"A35A63F5343EBE9EF8167BCB48AD122E"),
	(X"FFFFFFFFFFFFFFE00000000000000000", X"00000000000000000000000000000000", X"FD8687F0757A210E9FDF181204C30863"),
	(X"FFFFFFFFFFFFFFF00000000000000000", X"00000000000000000000000000000000", X"7A181E84BD5457D26A88FBAE96018FB0"),
	(X"FFFFFFFFFFFFFFF80000000000000000", X"00000000000000000000000000000000", X"653317B9362B6F9B9E1A580E68D494B5"),
	(X"FFFFFFFFFFFFFFFC0000000000000000", X"00000000000000000000000000000000", X"995C9DC0B689F03C45867B5FAA5C18D1"),
	(X"FFFFFFFFFFFFFFFE0000000000000000", X"00000000000000000000000000000000", X"77A4D96D56DDA398B9AABECFC75729FD"),
	(X"FFFFFFFFFFFFFFFF0000000000000000", X"00000000000000000000000000000000", X"84BE19E053635F09F2665E7BAE85B42D"),
	(X"FFFFFFFFFFFFFFFF8000000000000000", X"00000000000000000000000000000000", X"32CD652842926AEA4AA6137BB2BE2B5E"),
	(X"FFFFFFFFFFFFFFFFC000000000000000", X"00000000000000000000000000000000", X"493D4A4F38EBB337D10AA84E9171A554"),
	(X"FFFFFFFFFFFFFFFFE000000000000000", X"00000000000000000000000000000000", X"D9BFF7FF454B0EC5A4A2A69566E2CB84"),
	(X"FFFFFFFFFFFFFFFFF000000000000000", X"00000000000000000000000000000000", X"3535D565ACE3F31EB249BA2CC6765D7A"),
	(X"FFFFFFFFFFFFFFFFF800000000000000", X"00000000000000000000000000000000", X"F60E91FC3269EECF3231C6E9945697C6"),
	(X"FFFFFFFFFFFFFFFFFC00000000000000", X"00000000000000000000000000000000", X"AB69CFADF51F8E604D9CC37182F6635A"),
	(X"FFFFFFFFFFFFFFFFFE00000000000000", X"00000000000000000000000000000000", X"7866373F24A0B6ED56E0D96FCDAFB877"),
	(X"FFFFFFFFFFFFFFFFFF00000000000000", X"00000000000000000000000000000000", X"1EA448C2AAC954F5D812E9D78494446A"),
	(X"FFFFFFFFFFFFFFFFFF80000000000000", X"00000000000000000000000000000000", X"ACC5599DD8AC02239A0FEF4A36DD1668"),
	(X"FFFFFFFFFFFFFFFFFFC0000000000000", X"00000000000000000000000000000000", X"D8764468BB103828CF7E1473CE895073"),
	(X"FFFFFFFFFFFFFFFFFFE0000000000000", X"00000000000000000000000000000000", X"1B0D02893683B9F180458E4AA6B73982"),
	(X"FFFFFFFFFFFFFFFFFFF0000000000000", X"00000000000000000000000000000000", X"96D9B017D302DF410A937DCDB8BB6E43"),
	(X"FFFFFFFFFFFFFFFFFFF8000000000000", X"00000000000000000000000000000000", X"EF1623CC44313CFF440B1594A7E21CC6"),
	(X"FFFFFFFFFFFFFFFFFFFC000000000000", X"00000000000000000000000000000000", X"284CA2FA35807B8B0AE4D19E11D7DBD7"),
	(X"FFFFFFFFFFFFFFFFFFFE000000000000", X"00000000000000000000000000000000", X"F2E976875755F9401D54F36E2A23A594"),
	(X"FFFFFFFFFFFFFFFFFFFF000000000000", X"00000000000000000000000000000000", X"EC198A18E10E532403B7E20887C8DD80"),
	(X"FFFFFFFFFFFFFFFFFFFF800000000000", X"00000000000000000000000000000000", X"545D50EBD919E4A6949D96AD47E46A80"),
	(X"FFFFFFFFFFFFFFFFFFFFC00000000000", X"00000000000000000000000000000000", X"DBDFB527060E0A71009C7BB0C68F1D44"),
	(X"FFFFFFFFFFFFFFFFFFFFE00000000000", X"00000000000000000000000000000000", X"9CFA1322EA33DA2173A024F2FF0D896D"),
	(X"FFFFFFFFFFFFFFFFFFFFF00000000000", X"00000000000000000000000000000000", X"8785B1A75B0F3BD958DCD0E29318C521"),
	(X"FFFFFFFFFFFFFFFFFFFFF80000000000", X"00000000000000000000000000000000", X"38F67B9E98E4A97B6DF030A9FCDD0104"),
	(X"FFFFFFFFFFFFFFFFFFFFFC0000000000", X"00000000000000000000000000000000", X"192AFFFB2C880E82B05926D0FC6C448B"),
	(X"FFFFFFFFFFFFFFFFFFFFFE0000000000", X"00000000000000000000000000000000", X"6A7980CE7B105CF530952D74DAAF798C"),
	(X"FFFFFFFFFFFFFFFFFFFFFF0000000000", X"00000000000000000000000000000000", X"EA3695E1351B9D6858BD958CF513EF6C"),
	(X"FFFFFFFFFFFFFFFFFFFFFF8000000000", X"00000000000000000000000000000000", X"6DA0490BA0BA0343B935681D2CCE5BA1"),
	(X"FFFFFFFFFFFFFFFFFFFFFFC000000000", X"00000000000000000000000000000000", X"F0EA23AF08534011C60009AB29ADA2F1"),
	(X"FFFFFFFFFFFFFFFFFFFFFFE000000000", X"00000000000000000000000000000000", X"FF13806CF19CC38721554D7C0FCDCD4B"),
	(X"FFFFFFFFFFFFFFFFFFFFFFF000000000", X"00000000000000000000000000000000", X"6838AF1F4F69BAE9D85DD188DCDF0688"),
	(X"FFFFFFFFFFFFFFFFFFFFFFF800000000", X"00000000000000000000000000000000", X"36CF44C92D550BFB1ED28EF583DDF5D7"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFC00000000", X"00000000000000000000000000000000", X"D06E3195B5376F109D5C4EC6C5D62CED"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFE00000000", X"00000000000000000000000000000000", X"C440DE014D3D610707279B13242A5C36"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFF00000000", X"00000000000000000000000000000000", X"F0C5C6FFA5E0BD3A94C88F6B6F7C16B9"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFF80000000", X"00000000000000000000000000000000", X"3E40C3901CD7EFFC22BFFC35DEE0B4D9"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000", X"00000000000000000000000000000000", X"B63305C72BEDFAB97382C406D0C49BC6"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000", X"00000000000000000000000000000000", X"36BBAAB22A6BD4925A99A2B408D2DBAE"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000", X"00000000000000000000000000000000", X"307C5B8FCD0533AB98BC51E27A6CE461"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000", X"00000000000000000000000000000000", X"829C04FF4C07513C0B3EF05C03E337B5"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000", X"00000000000000000000000000000000", X"F17AF0E895DDA5EB98EFC68066E84C54"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000", X"00000000000000000000000000000000", X"277167F3812AFFF1FFACB4A934379FC3"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000", X"00000000000000000000000000000000", X"2CB1DC3A9C72972E425AE2EF3EB597CD"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000", X"00000000000000000000000000000000", X"36AEAA3A213E968D4B5B679D3A2C97FE"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000", X"00000000000000000000000000000000", X"9241DACA4FDD034A82372DB50E1A0F3F"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000", X"00000000000000000000000000000000", X"C14574D9CD00CF2B5A7F77E53CD57885"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000", X"00000000000000000000000000000000", X"793DE39236570ABA83AB9B737CB521C9"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000", X"00000000000000000000000000000000", X"16591C0F27D60E29B85A96C33861A7EF"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000", X"00000000000000000000000000000000", X"44FB5C4D4F5CB79BE5C174A3B1C97348"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000", X"00000000000000000000000000000000", X"674D2B61633D162BE59DDE04222F4740"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000", X"00000000000000000000000000000000", X"B4750FF263A65E1F9E924CCFD98F3E37"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000", X"00000000000000000000000000000000", X"62D0662D6EAEDDEDEBAE7F7EA3A4F6B6"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000", X"00000000000000000000000000000000", X"70C46BB30692BE657F7EAA93EBAD9897"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000", X"00000000000000000000000000000000", X"323994CFB9DA285A5D9642E1759B224A"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000", X"00000000000000000000000000000000", X"1DBF57877B7B17385C85D0B54851E371"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800", X"00000000000000000000000000000000", X"DFA5C097CDC1532AC071D57B1D28D1BD"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00", X"00000000000000000000000000000000", X"3A0C53FA37311FC10BD2A9981F513174"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00", X"00000000000000000000000000000000", X"BA4F970C0A25C41814BDAE2E506BE3B4"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00", X"00000000000000000000000000000000", X"2DCE3ACB727CD13CCD76D425EA56E4F6"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80", X"00000000000000000000000000000000", X"5160474D504B9B3EEFB68D35F245F4B3"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0", X"00000000000000000000000000000000", X"41A8A947766635DEC37553D9A6C0CBB7"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0", X"00000000000000000000000000000000", X"25D6CFE6881F2BF497DD14CD4DDF445B"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0", X"00000000000000000000000000000000", X"41C78C135ED9E98C096640647265DA1E"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8", X"00000000000000000000000000000000", X"5A4D404D8917E353E92A21072C3B2305"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC", X"00000000000000000000000000000000", X"02BC96846B3FDC71643F384CD3CC3EAF"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE", X"00000000000000000000000000000000", X"9BA4A9143F4E5D4048521C4F8877D88E"),
	(X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF", X"00000000000000000000000000000000", X"A1F6258C877D5FCD8964484538BFC92C")
    );
end package aes128Test;
